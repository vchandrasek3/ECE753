module TSC_16bit (f, g, x0, x1, y0, y1);

output f, g;

input [15:0] x0, x1, y0, y1;
//wire [29:0] a, b; 

wire [31:0] a, b;

/*
//Level 1
TSC T[15:0] (.f (f1[15:0]), .g (g1[15:0]), .x0 (x0[15:0]), .x1 (x1[15:0]), .y0 (y0[15:0]), .y1 (y1[15:0]) ); 

//Level 2
TSC L1 (.f (f2[0]), .g (g2[0]), .x0 (f1[0]), .y0 (g1[0]), .x1 (f1[1]), .y1 (g1[1]) );
TSC L2 (.f (f2[1]), .g (g2[1]), .x0 (f1[2]), .y0 (g1[2]), .x1 (f1[3]), .y1 (g1[3]) );
TSC L3 (.f (f2[2]), .g (g2[2]), .x0 (f1[4]), .y0 (g1[4]), .x1 (f1[5]), .y1 (g1[5]) );
TSC L4 (.f (f2[3]), .g (g2[3]), .x0 (f1[6]), .y0 (g1[6]), .x1 (f1[7]), .y1 (g1[7]) );
TSC L5 (.f (f2[4]), .g (g2[4]), .x0 (f1[8]), .y0 (g1[8]), .x1 (f1[9]), .y1 (g1[9]) );
TSC L6 (.f (f2[5]), .g (g2[5]), .x0 (f1[10]), .y0 (g1[10]), .x1 (f1[11]), .y1 (g1[11]) );
TSC L7 (.f (f2[6]), .g (g2[6]), .x0 (f1[12]), .y0 (g1[12]), .x1 (f1[13]), .y1 (g1[13]) );
TSC L8 (.f (f2[7]), .g (g2[7]), .x0 (f1[14]), .y0 (g1[14]), .x1 (f1[15]), .y1 (g1[15]) );

//Level 3
TSC M1 (.f (f3[0]), .g (g3[0]), .x0 (f2[0]), .y0 (g2[0]), .x1 (f2[1]), .y1 (g2[1]) );
TSC M2 (.f (f3[1]), .g (g3[1]), .x0 (f2[2]), .y0 (g2[2]), .x1 (f2[3]), .y1 (g2[3]) );
TSC M3 (.f (f3[2]), .g (g3[2]), .x0 (f2[4]), .y0 (g2[4]), .x1 (f2[5]), .y1 (g2[5]) );
TSC M4 (.f (f3[3]), .g (g3[3]), .x0 (f2[6]), .y0 (g2[6]), .x1 (f2[7]), .y1 (g2[7]) );

//Level 4
TSC N1 (.f (f4[0]), .g (g4[0]), .x0 (f3[0]), .y0 (g3[0]), .x1 (f3[1]), .y1 (g3[1]) );
TSC N2 (.f (f4[1]), .g (g4[1]), .x0 (f3[2]), .y0 (g3[2]), .x1 (f3[3]), .y1 (g3[3]) );

//Level 5 (Final)
TSC O1 (.f (f), .g (g), .x0 (f4[0]), .y0 (g4[0]), .x1 (f4[1]), .y1 (g4[1]) );
*/

TSC T00 (.f (a[0]), .g (b[0]), .x0 (x0[0]), .y0 (y0[0]), .x1 (x1[0]), .y1 (y1[0]) );
TSC T01 (.f (a[1]), .g (b[1]), .x0 (x0[1]), .y0 (y0[1]), .x1 (x1[1]), .y1 (y1[1]) );
TSC T02 (.f (a[2]), .g (b[2]), .x0 (a[0]), .y0 (b[0]), .x1 (a[1]), .y1 (b[1]) );
TSC T03 (.f (a[3]), .g (b[3]), .x0 (x0[2]), .y0 (y0[2]), .x1 (x1[2]), .y1 (y1[2]) );
TSC T04 (.f (a[4]), .g (b[4]), .x0 (a[2]), .y0 (b[2]), .x1 (a[3]), .y1 (b[3]) );
TSC T05 (.f (a[5]), .g (b[5]), .x0 (x0[3]), .y0 (y0[3]), .x1 (x1[3]), .y1 (y1[3]) );
TSC T06 (.f (a[6]), .g (b[6]), .x0 (a[4]), .y0 (b[4]), .x1 (a[5]), .y1 (b[5]) );
TSC T07 (.f (a[7]), .g (b[7]), .x0 (x0[4]), .y0 (y0[4]), .x1 (x1[4]), .y1 (y1[4]) );
TSC T08 (.f (a[8]), .g (b[8]), .x0 (a[6]), .y0 (b[6]), .x1 (a[7]), .y1 (b[7]) );
TSC T09 (.f (a[9]), .g (b[9]), .x0 (x0[5]), .y0 (y0[5]), .x1 (x1[5]), .y1 (y1[5]) );
TSC T10 (.f (a[10]), .g (b[10]), .x0 (a[8]), .y0 (b[8]), .x1 (a[9]), .y1 (b[9]) );
TSC T11 (.f (a[11]), .g (b[11]), .x0 (x0[6]), .y0 (y0[6]), .x1 (x1[6]), .y1 (y1[6]) );
TSC T12 (.f (a[12]), .g (b[12]), .x0 (a[10]), .y0 (b[10]), .x1 (a[11]), .y1 (b[11]) );
TSC T13 (.f (a[13]), .g (b[13]), .x0 (x0[7]), .y0 (y0[7]), .x1 (x1[7]), .y1 (y1[7]) );
TSC T14 (.f (a[14]), .g (b[14]), .x0 (a[12]), .y0 (b[12]), .x1 (a[13]), .y1 (b[13]) );
TSC T15 (.f (a[15]), .g (b[15]), .x0 (x0[8]), .y0 (y0[8]), .x1 (x1[8]), .y1 (y1[8]) );
TSC T16 (.f (a[16]), .g (b[16]), .x0 (a[14]), .y0 (b[14]), .x1 (a[15]), .y1 (b[15]) );
TSC T17 (.f (a[17]), .g (b[17]), .x0 (x0[9]), .y0 (y0[9]), .x1 (x1[9]), .y1 (y1[9]) );
TSC T18 (.f (a[18]), .g (b[18]), .x0 (a[16]), .y0 (b[16]), .x1 (a[17]), .y1 (b[17]) );
TSC T19 (.f (a[19]), .g (b[19]), .x0 (x0[10]), .y0 (y0[10]), .x1 (x1[10]), .y1 (y1[10]) );
TSC T20 (.f (a[20]), .g (b[20]), .x0 (a[18]), .y0 (b[18]), .x1 (a[19]), .y1 (b[19]) );
TSC T21 (.f (a[21]), .g (b[21]), .x0 (x0[11]), .y0 (y0[11]), .x1 (x1[11]), .y1 (y1[11]) );
TSC T22 (.f (a[22]), .g (b[22]), .x0 (a[20]), .y0 (b[20]), .x1 (a[21]), .y1 (b[21]) );
TSC T23 (.f (a[23]), .g (b[23]), .x0 (x0[12]), .y0 (y0[12]), .x1 (x1[12]), .y1 (y1[12]) );
TSC T24 (.f (a[24]), .g (b[24]), .x0 (a[22]), .y0 (b[22]), .x1 (a[23]), .y1 (b[23]) );
TSC T25 (.f (a[25]), .g (b[25]), .x0 (x0[13]), .y0 (y0[13]), .x1 (x1[13]), .y1 (y1[13]) );
TSC T26 (.f (a[26]), .g (b[26]), .x0 (a[24]), .y0 (b[24]), .x1 (a[25]), .y1 (b[25]) );
TSC T27 (.f (a[27]), .g (b[27]), .x0 (x0[14]), .y0 (y0[14]), .x1 (x1[14]), .y1 (y1[14]) );
TSC T28 (.f (a[28]), .g (b[28]), .x0 (a[26]), .y0 (b[26]), .x1 (a[27]), .y1 (b[27]) );
TSC T29 (.f (a[29]), .g (b[29]), .x0 (x0[15]), .y0 (y0[15]), .x1 (x1[15]), .y1 (y1[15]) );
//TSC T30 (.f (f), .g (g), .x0 (a[28]), .y0 (b[28]), .x1 (a[29]), .y1 (b[29]) );
TSC T30 (.f (a[30]), .g (b[30]), .x0 (a[28]), .y0 (b[28]), .x1 (a[29]), .y1 (b[29]) );
TSC T31 (.f (a[31]), .g (b[31]), .x0 (x0[0]), .y0 (y0[0]), .x1 (x1[0]), .y1 (y1[0]) );
TSC T32 (.f (f), .g (g), .x0 (a[30]), .y0 (b[30]), .x1 (a[31]), .y1 (b[31]) );



endmodule
