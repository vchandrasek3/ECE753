module TSC_16bit (f, g, x0, x1, y0, y1);

output f, g;

input [15:0] x0, x1, y0, y1;
wire [15:0] f1, g1;
wire [7:0] f2, g2;
wire [3:0] f3, g3;
wire [1:0] f4, g4;

//Level 1
TSC T[15:0] (.f (f1[15:0]), .g (g1[15:0]), .x0 (x0[15:0]), .x1 (x1[15:0]), .y0 (y0[15:0]), .y1 (y1[15:0]) ); 

//Level 2
TSC L1 (.f (f2[0]), .g (g2[0]), .x0 (f1[0]), .y0 (g1[0]), .x1 (f1[1]), .y1 (g1[1]) );
TSC L2 (.f (f2[1]), .g (g2[1]), .x0 (f1[2]), .y0 (g1[2]), .x1 (f1[3]), .y1 (g1[3]) );
TSC L3 (.f (f2[2]), .g (g2[2]), .x0 (f1[4]), .y0 (g1[4]), .x1 (f1[5]), .y1 (g1[5]) );
TSC L4 (.f (f2[3]), .g (g2[3]), .x0 (f1[6]), .y0 (g1[6]), .x1 (f1[7]), .y1 (g1[7]) );
TSC L5 (.f (f2[4]), .g (g2[4]), .x0 (f1[8]), .y0 (g1[8]), .x1 (f1[9]), .y1 (g1[9]) );
TSC L6 (.f (f2[5]), .g (g2[5]), .x0 (f1[10]), .y0 (g1[10]), .x1 (f1[11]), .y1 (g1[11]) );
TSC L7 (.f (f2[6]), .g (g2[6]), .x0 (f1[12]), .y0 (g1[12]), .x1 (f1[13]), .y1 (g1[13]) );
TSC L8 (.f (f2[7]), .g (g2[7]), .x0 (f1[14]), .y0 (g1[14]), .x1 (f1[15]), .y1 (g1[15]) );

//Level 3
TSC M1 (.f (f3[0]), .g (g3[0]), .x0 (f2[0]), .y0 (g2[0]), .x1 (f2[1]), .y1 (g2[1]) );
TSC M2 (.f (f3[1]), .g (g3[1]), .x0 (f2[2]), .y0 (g2[2]), .x1 (f2[3]), .y1 (g2[3]) );
TSC M3 (.f (f3[2]), .g (g3[2]), .x0 (f2[4]), .y0 (g2[4]), .x1 (f2[5]), .y1 (g2[5]) );
TSC M4 (.f (f3[3]), .g (g3[3]), .x0 (f2[6]), .y0 (g2[6]), .x1 (f2[7]), .y1 (g2[7]) );

//Level 4
TSC N1 (.f (f4[0]), .g (g4[0]), .x0 (f3[0]), .y0 (g3[0]), .x1 (f3[1]), .y1 (g3[1]) );
TSC N2 (.f (f4[1]), .g (g4[1]), .x0 (f3[2]), .y0 (g3[2]), .x1 (f3[3]), .y1 (g3[3]) );

//Level 5 (Final)
TSC O1 (.f (f), .g (g), .x0 (f4[0]), .y0 (g4[0]), .x1 (f4[1]), .y1 (g4[1]) );



endmodule
