module TSC_Reconfig_tb();

wire [15:0] final_x, final_y;
reg [15:0] x0, x1, y0, y1;

TSC_Reconfig U0 (.final_x(final_x), .final_y(final_y), .x0(x0), .y0(y0), .x1(x1), .y1(y1));

initial begin
//0000
x0 = 16'b0000000000000000;
y0 = 16'b0000000000000000;
x1 = 16'b0000000000000000;
y1 = 16'b0000000000000000;

//0001
#10
x0 = 16'b0000000000000000;
y0 = 16'b0000000000000000;
x1 = 16'b0000000000000000;
y1 = 16'b1111111111111111;

//0010
#10
x0 = 16'b0000000000000000;
y0 = 16'b0000000000000000;
x1 = 16'b1111111111111111;
y1 = 16'b0000000000000000;

//0011
#10
x0 = 16'b0000000000000000;
y0 = 16'b0000000000000000;
x1 = 16'b1111111111111111;
y1 = 16'b1111111111111111;

//0100
#10
x0 = 16'b0000000000000000;
y0 = 16'b1111111111111111;
x1 = 16'b0000000000000000;
y1 = 16'b0000000000000000;

//0101 CODEWORD
#10
x0 = 16'b0000000000000000;
y0 = 16'b1111111111111111;
x1 = 16'b0000000000000000;
y1 = 16'b1111111111111111;

//0110 CODEWORD
#10
x0 = 16'b0000000000000000;
y0 = 16'b1111111111111111;
x1 = 16'b1111111111111111;
y1 = 16'b0000000000000000;

//0111 
#10
x0 = 16'b0000000000000000;
y0 = 16'b1111111111111111;
x1 = 16'b1111111111111111;
y1 = 16'b1111111111111111;

//1000
#10
x0 = 16'b1111111111111111;
y0 = 16'b0000000000000000;
x1 = 16'b0000000000000000;
y1 = 16'b0000000000000000;

//1001 CODEWORD
#10
x0 = 16'b1111111111111111;
y0 = 16'b0000000000000000;
x1 = 16'b0000000000000000;
y1 = 16'b1111111111111111;

//1010 CODEWORD
#10
x0 = 16'b1111111111111111;
y0 = 16'b0000000000000000;
x1 = 16'b1111111111111111;
y1 = 16'b0000000000000000;

//1011
#10
x0 = 16'b1111111111111111;
y0 = 16'b0000000000000000;
x1 = 16'b1111111111111111;
y1 = 16'b1111111111111111;

//1100
#10
x0 = 16'b1111111111111111;
y0 = 16'b1111111111111111;
x1 = 16'b0000000000000000;
y1 = 16'b0000000000000000;

//1101
#10
x0 = 16'b1111111111111111;
y0 = 16'b1111111111111111;
x1 = 16'b0000000000000000;
y1 = 16'b1111111111111111;

//1110
#10
x0 = 16'b1111111111111111;
y0 = 16'b1111111111111111;
x1 = 16'b1111111111111111;
y1 = 16'b0000000000000000;

//1111
#10
x0 = 16'b1111111111111111;
y0 = 16'b1111111111111111;
x1 = 16'b1111111111111111;
y1 = 16'b1111111111111111;

end

initial  begin
$display("\tTIME, \tx0, \ty0, \tx1, \ty1, \tfinal_x, \tfinal_y, \tlogic_en, \tf, \tg"); 
$monitor("%d,\t%b,\t%b,\t%b,\t%b, \t%b,\t%b, \t%b, \t%b, \t%b",$time, x0, y0, x1, y1, final_x, final_y, U0.logic_en, U0.DUT1.f, U0.DUT1.g); 
end 

endmodule
